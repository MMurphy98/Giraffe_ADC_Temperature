module Giraffe_FSM #(
    parameters
) (
    ports
);

endmodule